module ctrl
(

);

endmodule