`define datawidth 30