`define datawidth 14